** sch_path: /home/tare/ITI_Analog/ITI_Labs/Lab4/Design/Lab04.sch
**.subckt Lab04
V1 VSIG GND AC 1
I0 VDD VOUT 10u
V2 VDD GND 1.8
RSIG VIN VSIG 2meg m=1
XM0 GND VIN VOUT VOUT pmos_3p3 L=1u W=20u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
C1 VOUT GND 2p m=1
**** begin user architecture code

.include /home/tare/pdk/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/tare/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include sim_script.sim


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
