** sch_path: /home/tare/Desktop/ITI_Analog/ITI_Labs/Lab5/Design/Lab5.sch
**.subckt Lab5
XM0 net1 net1 GND GND nmos_3p3 L=1.42u W=14.58u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
VDD VDD GND 1.8
IB1 VDD net1 10u
VGMIS net2 net1 0
VOUT VOUT GND 0.9
RB net7 net4 20k m=1
XM1 VOUT net2 GND GND nmos_3p3 L=1.42u W=2*14.58u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
IB2 VDD net7 10u
XM2 net3 net4 GND GND nmos_3p3 L=1.42u W=14.58u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM3 VDS3 net6 GND GND nmos_3p3 L=1.42u W=2*14.58u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM4 net4 net7 net3 GND nmos_3p3 L=1.42u W=14.58u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM5 VOUT net5 VDS3 GND nmos_3p3 L=1.42u W=2*14.58u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
VGMIS1 net6 net4 0
VGMIS2 net5 net7 0
**** begin user architecture code


.include sim_script.sim



.include /home/tare/pdk/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/tare/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
