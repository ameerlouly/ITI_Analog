** sch_path: /home/tare/ITI_Analog/ITI_Labs/Lab1/RC/Design/RC.sch
**.subckt RC
C1 VOUT GND 1p m=1
R1 VOUT VIN 1k m=1
V2 VIN GND DC 0 AC 1
**** begin user architecture code


.control
ac dec 10 1 10G
save all
meas ac MAX_GAIN MAX vmag(vout) from=1 to=10G
meas ac BW when vmag(vout)=0.707 fall = 1
write rc_ckt_ac.raw
set appendwrite
touch ac_results.txt
print MAX_GAIN BW > ac_results.txt
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
