** sch_path: /home/tare/ITI_Analog/Lab2/Design/Lab02_DC.sch
**.subckt Lab02_DC
VIN VIN GND DC 0 AC 1
V2 VDD GND 2.5
R3 VDD VOUT 100k m=1
XM1 VOUT VIN GND GND nmos_3p3 L=2u W=9.76u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
**** begin user architecture code

.include /home/tare/pdk/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/tare/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.control
save all
+ @m.xm1.m0[id]
+ @m.xm1.m0[gm]
+ @m.xm1.m0[gds]
+ @m.xm1.m0[vgs]
+ @m.xm1.m0[vds]
dc VIN 0 2.5 10m
remzerovec
write Lab02_DC.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
